----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    09:19:25 10/20/2017 
-- Design Name: 
-- Module Name:    DataMemory - tbDataMemory 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.all;
use IEEE.std_logic_unsigned.all;


entity DataMemory is
    Port ( cRD : in  STD_LOGIC_VECTOR (31 downto 0);
           AluResult : in  STD_LOGIC_VECTOR (31 downto 0);
           WRENMEM : in  STD_LOGIC;
			  Reset : in STD_LOGIC;
           DataMem : out  STD_LOGIC_VECTOR (31 downto 0));
end DataMemory;

architecture Behavioral of DataMemory is

type reg is array (0 to 519) of std_logic_vector (31 downto 0);
signal myReg : reg := (others => x"00000000");

begin

process(cRD,AluResult,Reset,WRENMEM) begin
	if (Reset = '1') then
		myReg <= (others => x"00000000");
	else 
		if (WRENMEM = '1') then
			myReg(conv_integer(AluResult)) <= cRD;
		end if;
		if(520>AluResult) then
			DataMem <= myReg(conv_integer(AluResult));
		end if;
	end if;
end process;



end Behavioral;
