----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    10:51:25 10/20/2017 
-- Design Name: 
-- Module Name:    MuxRF - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity MuxRF is
    Port ( Rd : in  STD_LOGIC_VECTOR (5 downto 0);
           O7 : in  STD_LOGIC_VECTOR (5 downto 0);
           RFDEST : in  STD_LOGIC;
           nRD : out  STD_LOGIC_VECTOR (5 downto 0));
end MuxRF;

architecture Behavioral of MuxRF is
signal nRD_Aux : STD_LOGIC_VECTOR (5 downto 0) := "000000";
begin
	process (Rd,O7,RFDEST) begin
		
		case (RFDEST) is 
		when '0' => 
		nRD <= Rd;
		when '1' =>
		nRD <= O7;
		when others => 
		nRD <= Rd;
	end case;
	
end process;


end Behavioral;


