----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    16:37:34 09/26/2017 
-- Design Name: 
-- Module Name:    IM - Arqim 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

use ieee.std_logic_unsigned.all;
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity IM is
    Port ( Address : in  STD_LOGIC_VECTOR (31 downto 0);
           Reset : in  STD_LOGIC;
           Instruction : out  STD_LOGIC_VECTOR (31 downto 0));
end IM;

architecture Arqim of IM is

type rom_type is array (63 downto 0) of std_logic_vector (31 downto 0);
signal ROM : rom_type := (	"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"00000000000000000000000000000000", "00000000000000000000000000000000",
									"10010110000100000000000000001010", "10111000000100000010000000000011",
									"01111111111111111111111111101111", "10110110000100000010000000000010",
									"10010100000100000000000000010011", "10000001110000111110000000000001",
									"00000001000000000000000000000000", "00010000101111111111111111110110",
									"10101010000100000000000000000011", "10000110000001010110000000000001",
									"10100110000100000000000000001001", "00000001000000000000000000000000",
									"01111111111111111111111111101100", "10110100000100000000000000011011",
									"10110010000100000000000000010011", "00000001000000000000000000000000",
									"00010110100000000000000000001011", "10000000101001010100000000011100",
									"10101010000100000010000000000000", "10100110000100000010000000000001",
									"10010010000100000000000000010001", "10000001110000111110000000000001",
									"00000001000000000000000000000000", "00110000101111111111111111111001",
									"10100100000100000000000000000010", "10000100000001001010000000000001",
									"10100010000100000000000000000001", "10000010000001000100000000011001",
									"00000001000000000000000000000000", "00110110100000000000000000001000",
									"10000000101001001000000000011010", "10100100000100000010000000000000",
									"10100010000100000010000000000000", "00010000100000000000000000011110");

begin

    process (Reset,Address,rom)
    begin
        if (Reset='1') then
				Instruction <= "00000000000000000000000000000000";
		  else
            Instruction <= ROM(conv_integer(Address(5 downto 0)));  
        end if;
    end process;
end Arqim;

